module top(output led);
   assign led=1;
endmodule
